module dbi_tx_fsm 
#(

) (

);

endmodule