module axi4_fifo 
#(

) (

);

endmodule