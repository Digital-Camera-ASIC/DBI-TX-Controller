module dbi_tx_phy 
#(

) (

);

endmodule